module and_4bit(y,a,b,c,d);
input a,b,c,d;
output y;
assign y = a&b&c&d;
endmodule
